`include "constants.vh"
`default_nettype none
module alu_src_a_mux (
    
    );

endmodule

module alu_src_b_mux (

    );

endmodule

module mul_src_a_mux (

    );

endmodule

