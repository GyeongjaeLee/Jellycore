`include "constants.vh"
`default_nettype none
module prefix_sum(
    input wire  [`IQ_ENT_NUM-1:0]   request,
    output wire                     grant,
    output wire [`IQ_ENT_SEL-1:0]   selected_ent
    );

endmodule